`ifndef APB_IFS__SV
`define APB_IFS__SV 

interface apb_ifs;

endinterface

`endif
