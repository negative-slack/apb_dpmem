`ifndef APB_DPMEM_ENV__SV
`define APB_DPMEM_ENV__SV 

class apb_dpmem_env extends uvm_env;

  //////////////////////////////////////////////////////////////////////////////
  // Declaration of component utils to register with factory 
  //////////////////////////////////////////////////////////////////////////////
  `uvm_component_utils(apb_dpmem_env)

  //////////////////////////////////////////////////////////////////////////////
  // agent and scoreboard instance
  //////////////////////////////////////////////////////////////////////////////
  apb_dpmem_agent      apb_dpmem_agnt;
  apb_dpmem_ref_model  apb_dpmem_rm;
  apb_dpmem_scoreboard apb_dpmem_scb;

  ///////////////////////////////////////////////////////////////////////////////
  // Method name : new 
  // Description : constructor
  ///////////////////////////////////////////////////////////////////////////////
  function new(string name, uvm_component parent);
    super.new(name, parent);
  endfunction : new

  ///////////////////////////////////////////////////////////////////////////////
  // Method name : build-phase 
  // Description : construct the components such as.. agent, scoreboard 
  ///////////////////////////////////////////////////////////////////////////////
  function void build_phase(uvm_phase phase);
    super.build_phase(phase);
    apb_dpmem_agnt = mem_agent::type_id::create("apb_dpmem_agnt", this);
    apb_dpmem_scb  = mem_scoreboard::type_id::create("apb_dpmem_scb", this);
  endfunction : build_phase

  ///////////////////////////////////////////////////////////////////////////////
  // Method name : connect_phase 
  // Description : connect tlm ports ande exports (ex: analysis port/exports) 
  ///////////////////////////////////////////////////////////////////////////////
  function void connect_phase(uvm_phase phase);
    apb_dpmem_agnt.monitor.item_collected_port.connect(apb_dpmem_scb.item_collected_export);
  endfunction : connect_phase

endclass : mem_model_env

`endif
