`ifndef APV_IF_DV__SV
`define APV_IF_DV__SV 

class apb_if_dv extends apb_if;

endclass : apb_if_dv

`endif
