`ifndef APB_DPMEM_REF_MODEL_PKG__SV
`define APB_DPMEM_REF_MODEL_PKG__SV 

package apb_dpmem_ref_model_pkg;
  `include "uvm_macros.svh"
  import uvm_pkg::*;

  //////////////////////////////////////////////////////////
  // importing packages : agent, ref model
  /////////////////////////////////////////////////////////
  import apb_dpmem_agent_pkg::*;

  //////////////////////////////////////////////////////////
  // include ref model files 
  /////////////////////////////////////////////////////////
  `include "apb_dpmem_ref_model.sv"

endpackage

`endif

