`ifndef APB_DPMEM_AGENT__SV
`define APB_DPMEM_AGENT__SV 

class apb_dpmem_agent extends uvm_agent;

  ///////////////////////////////////////////////////////////////////////////////
  // Declaration of component utils 
  ///////////////////////////////////////////////////////////////////////////////
  `uvm_component_utils(apb_dpmem_agent)

  ///////////////////////////////////////////////////////////////////////////////
  // Method name : new 
  // Description : constructor
  ///////////////////////////////////////////////////////////////////////////////
  function new(string name, uvm_component parent);
    super.new(name, parent);
  endfunction : new

  ///////////////////////////////////////////////////////////////////////////////
  // Declaration of UVM components such as.. driver, sequencer, monitor 
  ///////////////////////////////////////////////////////////////////////////////
  apb_dpmem_sequencer sequencer;
  apb_dpmem_driver    driver;
  apb_dpmem_monitor   monitor;

  ///////////////////////////////////////////////////////////////////////////////
  // Method name : build-phase 
  // Description : construct the components such as.. driver, sequencer, monitor
  ///////////////////////////////////////////////////////////////////////////////
  function void build_phase(uvm_phase phase);
    super.build_phase(phase);
    sequencer = apb_dpmem_sequencer::type_id::create("sequencer", this);
    driver = apb_dpmem_driver::type_id::create("driver", this);
    monitor = apb_dpmem_monitor::type_id::create("monitor", this);
  endfunction : build_phase

  ///////////////////////////////////////////////////////////////////////////////
  // Method name : connect_phase 
  // Description : connect the export of the sequence to the port of the driver 
  //               that's how the transactions are sent !  
  ///////////////////////////////////////////////////////////////////////////////
  function void connect_phase(uvm_phase phase);
    driver.seq_item_port.connect(sequencer.seq_item_export);
  endfunction : connect_phase

endclass : apb_dpmem_agent

`endif
